`ifndef PB_UVC_PKG
`define PB_UVC_PKG

`inculde "pb_interface.sv"

package pb_uvc_pkg;

`include "uvm_macros.svh"
import uvm_pkg::*;

`include "pb_common.sv"
`include "pb_agent_cfg.sv"
`include "pb_item.sv"
`include "pb_monitor.sv"
`include "pb_agent.sv"
`include "pb_env.sv"

endpackage : pb_uvc_pkg

`endif // PB_UVC_pkg