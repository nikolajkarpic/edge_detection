`ifndef ITEM
`define ITEM

class item extends uvm_sequence_item;

    //fields

    // registration macros
    `uvm_component_utils_begin(item)
        //field registration
    `uvm_component_utils_end

endclass : item

`endif // item