`ifndef UVC_PKG
`define UVC_PKG

`inculde "interface.sv"

package uvc_pkg;

`include "uvm_macros.svh"
import uvm_pkg::*;

// `include "common.sv"
`include "agent_cfg.sv"
`include "item.sv"
`include "driver.sv"
`include "sequencer.sv"
`include "monitor.sv"
//`include "cov.sv"
`include "agent.sv"
`include "env.sv"
`include "seq_lib.sv"

endpackage : uvc_pkg

`endif // UVC_pkg