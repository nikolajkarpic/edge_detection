`ifndef COMMON
`define COMMON



`endif // COMMON