`ifndef END_COMMON
`define END_COMMON

typedef enum {IN_DAT, OUT_DAT, START, DONE} end_trans_type;

bit [7:0] img1 [10000] = '{
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01111011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"01111011",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"11111111",
"01111011",
"11111111",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"01111011",
"01111011",
"01111011",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"01111011",
"01111011",
"01111011",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"01111011",
"01111011",
"01111011",
"11111111",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"11111111",
"01111011",
"01111011",
"01111011",
"11111111",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"11111111",
"11111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"11111111",
"11111111",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"11111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"11111111",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"11111111",
"11111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"11111111",
"11111111",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"11111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"11111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"11111111",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"11111111",
"01111011",
"01111011",
"01111011",
"01111011",
"11111111",
"11111111",
"11111111",
"01111011",
"01111011",
"01111011",
"01111011",
"11111111",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"11111111",
"11111111",
"01111011",
"01111011",
"01111011",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"01111011",
"01111011",
"01111011",
"11111111",
"11111111",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"11111111",
"11111111",
"01111011",
"01111011",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"01111011",
"01111011",
"11111111",
"11111111",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"11111111",
"01111011",
"01111011",
"11111111",
"11111111",
"11111111",
"11111111",
"11001001",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"01111011",
"11111111",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11111111",
"11111111",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11111111",
"11111111",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11111111",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11111111",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"11001001",
"11001001",
"11001001",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"11001001",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01011011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01011011",
"01011011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111011",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111011",
"01111011",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111",
"01111111"
};

`endif // END_COMMON