`ifndef test_pkg
`define test_pkg

package test_pkg;

`include "uvm_macros.svh"
import uvm_pkg::*;

import addr_uvc_pkg::*;
import end_uvc_pkg::*;
import mem_uvc_pkg::*;
import pb_uvc_pkg::*;

import top_env_pkg::*;

//include sequences
`include "test_base.sv"
`include "test_img.sv"
// include tests

endpackage : test_pkg

`endif // test_pkg