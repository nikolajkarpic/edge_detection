`ifndef PB_COMMON
`define PB_COMMON

typedef enum {DAT,EN,SUM_OUT} pb_packet_type;

`endif // PB_COMMON