`ifndef ADDR_COMMON
`define ADDR_COMMON

typedef enum {CALC_CONV,CALC_ADDR,SHIFT} addr_packet_type;

`endif // ADDR_COMMON