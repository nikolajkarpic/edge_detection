`ifndef MEM_COMMON
`define MEM_COMMON

typedef enum {SHIFT,DAT_OUT,KERN_OUT} mem_packet_type;

`endif // MEM_COMMON