`ifndef INTERFACE
`define INTERFACE

interface intf(input CLK, input RST);

    `include "uvm_macros.svh"

    // signals

endinterface : intf

`endif // INTERFACE