`ifndef ADDR_COMMON
`define ADDR_COMMON

typedef enum {CALC_CONV,CALC_ADDR,SHIFTING} addr_packet_type;
typedef enum {ACTIVE,PASIVE} active_pasive;

`endif // ADDR_COMMON